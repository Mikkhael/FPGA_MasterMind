parameter ADDR_W = 4'd9;
parameter FONT_H = 3'd5;
parameter FONT_W = 3'd4;
parameter FONT_CHARS = 6'd44;
parameter FONT_LINEOFF = 7'd64;
parameter FONT_LINESHIFT = 3'd6;
parameter CHAR_0 = 1'd0;
parameter CHAR_1 = 1'd1;
parameter CHAR_2 = 2'd2;
parameter CHAR_3 = 2'd3;
parameter CHAR_4 = 3'd4;
parameter CHAR_5 = 3'd5;
parameter CHAR_6 = 3'd6;
parameter CHAR_7 = 3'd7;
parameter CHAR_8 = 4'd8;
parameter CHAR_9 = 4'd9;
parameter CHAR_A = 4'd10;
parameter CHAR_B = 4'd11;
parameter CHAR_C = 4'd12;
parameter CHAR_D = 4'd13;
parameter CHAR_E = 4'd14;
parameter CHAR_F = 4'd15;
parameter CHAR_G = 5'd16;
parameter CHAR_H = 5'd17;
parameter CHAR_I = 5'd18;
parameter CHAR_J = 5'd19;
parameter CHAR_K = 5'd20;
parameter CHAR_L = 5'd21;
parameter CHAR_M = 5'd22;
parameter CHAR_N = 5'd23;
parameter CHAR_O = 5'd24;
parameter CHAR_P = 5'd25;
parameter CHAR_Q = 5'd26;
parameter CHAR_R = 5'd27;
parameter CHAR_S = 5'd28;
parameter CHAR_T = 5'd29;
parameter CHAR_U = 5'd30;
parameter CHAR_V = 5'd31;
parameter CHAR_W = 6'd32;
parameter CHAR_X = 6'd33;
parameter CHAR_Y = 6'd34;
parameter CHAR_Z = 6'd35;
parameter CHAR_  = 6'd36;
parameter CHAR_QMark = 6'd37;
parameter CHAR_Hash = 6'd38;
parameter CHAR_Exclemation = 6'd39;
parameter CHAR_Colon = 6'd40;
parameter CHAR_LeftBracket = 6'd41;
parameter CHAR_ArrowR = 6'd42;
parameter CHAR_ArrowL = 6'd43;
parameter LSPRITE_MM_LEN = 2'd2;
parameter LSPRITE_Mind_LEN = 3'd4;
parameter LSPRITE_exit_LEN = 3'd4;
parameter LSPRITE_Enter_LEN = 2'd2;
parameter LSPRITE_MM = 6'd44;
parameter LSPRITE_Mind = 6'd46;
parameter LSPRITE_exit = 6'd50;
parameter LSPRITE_Enter = 6'd54;
parameter STR_TITLE_LEN = 4'd11;
parameter STR_PLAYVSCOMPUTER_LEN = 5'd16;
parameter STR_PLAYVSHUMAN_LEN = 4'd13;
parameter STR_PLAYVSRIVAL_LEN = 5'd25;
parameter STR_OPTIONS_LEN = 3'd7;
parameter STR_HIGHSCORES_LEN = 4'd10;
parameter STR_GUESS_LEN = 2'd2;
parameter STR_EXIT_LEN = 1'd1;
parameter STR_BACK_LEN = 4'd10;
parameter STR_YOUWIN_LEN = 4'd9;
parameter STR_GAMEOVER_LEN = 4'd12;
parameter STR_ENTERSECRET_LEN = 4'd13;
parameter STR_HINTSGREEN_LEN = 4'd13;
parameter STR_HINTSYELLOW_LEN = 4'd13;
parameter STR_GUESSER_LEN = 4'd13;
parameter STR_SETTER_LEN = 4'd12;
parameter STR_PINCOLORS_LEN = 4'd10;
parameter STR_PINSCOUNT_LEN = 4'd10;
parameter STR_GUESSES_LEN = 3'd7;
parameter STR_PIXELWIDTH_LEN = 4'd11;
parameter STR_PIXELHEIGHT_LEN = 4'd12;
parameter STR_PALETTE_LEN = 3'd7;
parameter logic [8:0] STR_TITLE [11] = '{44,45,10,28,29,14,27,46,47,48,49};
parameter logic [8:0] STR_PLAYVSCOMPUTER [16] = '{25,21,10,34,36,31,28,36,12,24,22,25,30,29,14,27};
parameter logic [8:0] STR_PLAYVSHUMAN [13] = '{25,21,10,34,36,31,28,36,17,30,22,10,23};
parameter logic [8:0] STR_PLAYVSRIVAL [25] = '{25,21,10,34,36,31,28,36,17,30,22,10,23,40,36,27,18,31,10,21,36,22,24,13,14};
parameter logic [8:0] STR_OPTIONS [7] = '{24,25,29,18,24,23,28};
parameter logic [8:0] STR_HIGHSCORES [10] = '{17,18,16,17,28,12,24,27,14,28};
parameter logic [8:0] STR_GUESS [2] = '{54,55};
parameter logic [8:0] STR_EXIT [1] = '{33};
parameter logic [8:0] STR_BACK [10] = '{43,43,36,11,10,12,20,36,43,43};
parameter logic [8:0] STR_YOUWIN [9] = '{34,24,30,36,32,18,23,39,39};
parameter logic [8:0] STR_GAMEOVER [12] = '{16,10,22,14,36,24,31,14,27,36,40,41};
parameter logic [8:0] STR_ENTERSECRET [13] = '{14,23,29,14,27,36,28,14,12,27,14,29,40};
parameter logic [8:0] STR_HINTSGREEN [13] = '{17,18,23,29,28,36,16,27,14,14,23,40,36};
parameter logic [8:0] STR_HINTSYELLOW [13] = '{17,18,23,29,28,36,34,14,21,21,24,32,40};
parameter logic [8:0] STR_GUESSER [13] = '{16,30,14,28,28,14,27,36,32,18,23,28,39};
parameter logic [8:0] STR_SETTER [12] = '{28,14,29,29,14,27,36,32,18,23,28,39};
parameter logic [8:0] STR_PINCOLORS [10] = '{25,18,23,36,12,24,21,24,27,28};
parameter logic [8:0] STR_PINSCOUNT [10] = '{25,18,23,28,36,12,24,30,23,29};
parameter logic [8:0] STR_GUESSES [7] = '{16,30,14,28,28,14,28};
parameter logic [8:0] STR_PIXELWIDTH [11] = '{25,18,33,14,21,36,32,18,13,29,17};
parameter logic [8:0] STR_PIXELHEIGHT [12] = '{25,18,33,14,21,36,17,14,18,16,17,29};
parameter logic [8:0] STR_PALETTE [7] = '{25,10,21,14,29,29,14};
parameter logic STR_MASK_TITLE [11] = '{1,0,0,0,0,0,0,1,1,1,0};
parameter logic STR_MASK_PLAYVSCOMPUTER [16] = '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_PLAYVSHUMAN [13] = '{0,0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_PLAYVSRIVAL [25] = '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_OPTIONS [7] = '{0,0,0,0,0,0,0};
parameter logic STR_MASK_HIGHSCORES [10] = '{0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_GUESS [2] = '{1,0};
parameter logic STR_MASK_EXIT [1] = '{0};
parameter logic STR_MASK_BACK [10] = '{0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_YOUWIN [9] = '{0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_GAMEOVER [12] = '{0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_ENTERSECRET [13] = '{0,0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_HINTSGREEN [13] = '{0,0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_HINTSYELLOW [13] = '{0,0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_GUESSER [13] = '{0,0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_SETTER [12] = '{0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_PINCOLORS [10] = '{0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_PINSCOUNT [10] = '{0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_GUESSES [7] = '{0,0,0,0,0,0,0};
parameter logic STR_MASK_PIXELWIDTH [11] = '{0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_PIXELHEIGHT [12] = '{0,0,0,0,0,0,0,0,0,0,0,0};
parameter logic STR_MASK_PALETTE [7] = '{0,0,0,0,0,0,0};
