parameter STR_TITLE_LEN = 12;
parameter logic [5:0] STR_TITLE [12] = '{36,37,10,28,29,14,27,36,37,18,23,13};
parameter STR_OPTS_LEN = 7;
parameter logic [5:0] STR_OPTS [7] = '{24,25,29,18,24,23,28};
parameter STR_TEST_LEN = 4;
parameter logic [5:0] STR_TEST [4] = '{29,14,28,29};
